module mult (
input i_x,
input i_y,
output [1:0] o_z
);

assign o_z = i_x * i_y;

endmodule
